`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: Maven Silicon -VIT Vellore
// Engineer: VLSI Design
// 
// Create Date: 26.06.2024 16:36:41
// Design Name: Instruction mux
// Module Name: msrv32_instruction_mux
// Project Name: RSIC -V 32I
// Target Devices: 
// Tool Versions: Achyut's Vivado
// Description: 
// RTL / design code
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module msrv32_instruction_mux(flush_in, ms_riscv32_mp_instr_in, opcode_out, funct3_out, funct7_out, rs1addr_out, rs2addr_out, rdaddr_out, csr_addr_out, instr_out);
input flush_in;
input [31:0] ms_riscv32_mp_instr_in;

output [6:0] opcode_out;
output [2:0] funct3_out;
output [6:0] funct7_out; 
output [4:0] rs1addr_out; 
output [4:0] rs2addr_out;
output [4:0] rdaddr_out;
output [11:0] csr_addr_out;
output [24:0]  instr_out;
wire [31:0] instr_mux;
assign  instr_mux = (flush_in)? 32'h00000013 : ms_riscv32_mp_instr_in;
assign opcode_out = instr_mux[6:0];
assign funct3_out = instr_mux[14:12];
assign funct7_out = instr_mux[31:25];
assign rs1addr_out = instr_mux[19:15];
assign rs2addr_out = instr_mux[24:20];
assign rdaddr_out = instr_mux[11:7];
assign csr_addr_out = instr_mux[31:20];
assign instr_out = instr_mux[31:7];
endmodule 
